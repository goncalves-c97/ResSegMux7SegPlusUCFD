----------------------------------------------------------------------------------
-- Company: Funda��o Engenheiro Salvador Arena 
--
-- Engineers: Carlos Adonias
--			  	  Carlos Gon�alves
--			 	  Gabriel Teixeira
-- 		 	  Johnny Messias
--
-- Teacher: Filippo Valiante
-- Create Date:    20:03:38 05/05/2023 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity FD_MUX is
end FD_MUX;

architecture Behavioral of FD_MUX is

begin


end Behavioral;

